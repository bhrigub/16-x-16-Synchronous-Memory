library verilog;
use verilog.vl_types.all;
entity tbm is
end tbm;
